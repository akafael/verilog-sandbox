/*
 * Very basic module
 *
 * @author Akafael
 */

module hello;
  initial 
    begin
      $display("Hello, World");
      $finish ;
    end
endmodule
